library ieee;
use ieee.std_logic_1164.all;

package core_pack is

  subtype dw_t is std_logic_vector(31 downto 0);

end package;
